module hf_compression ();

endmodule